`include "parameters.vh"

module display_ctrl(
    input clk,
    input rst,
    input [3:0] state,
    input [7:0] countdown,
    input [31:0] cycles,
    input [2:0] alu_op,
    input error_led,  // �������������LED�źţ�ά�Ȼ�������Чʱ������
    output reg [7:0] seg,
    output reg [3:0] an,
    output reg [7:0] led
);

    reg [1:0] scan_cnt; 
    reg [19:0] refresh_cnt; 

    reg [4:0] digit_0, digit_1, digit_2, digit_3; 
    reg [4:0] current_digit;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            digit_0 <= 5'h0F;
            digit_1 <= 5'h0F;
            digit_2 <= 5'h0F;
            digit_3 <= 5'h0F;
        end
        else begin
            
            digit_3 <= 5'h0F; digit_2 <= 5'h0F; digit_1 <= 5'h0F; digit_0 <= 5'h0F;

            case (state)
                `IDLE: begin
                    digit_3 <= 5'h01;  // I
                    digit_2 <= 5'h0D;  // d
                    digit_1 <= 5'h12;  // L
                    digit_0 <= 5'h0E;  // E
                end

                `INPUT_DIM, `INPUT_DATA, `FILL_ZEROS: begin
                    digit_3 <= 5'h01;  // I
                    digit_2 <= 5'h05;  // n
                    digit_1 <= 5'h10;  // P
                    digit_0 <= 5'h11;  // t
                end

                `COMPUTE: begin
                    // ��ʾ "CAL" + ��������
                    digit_3 <= 5'h0C;  // C
                    digit_2 <= 5'h0A;  // A
                    digit_1 <= 5'h12;  // L
                    // digit_0 ���� alu_op ��ʾ��������
                    // ����ͼƬҪ��0=T(CALT), 1=A(CALA), 2=b(CALb), 3=C(CALC), 4=J(CALJ)
                    case (alu_op)
                        3'd0: digit_0 <= 5'h14; // T
                        3'd1: digit_0 <= 5'h0A; // A
                        3'd2: digit_0 <= 5'h0B; // b (Сд)
                        3'd3: digit_0 <= 5'h0C; // C
                        3'd4: digit_0 <= 5'h15; // J
                        default: digit_0 <= 5'h0F; // F (��Ч����)
                    endcase
                end

                `DISPLAY_MODE: begin
                    
                    digit_3 <= 5'h0D;  // d
                    digit_2 <= 5'h01;  // I
                    digit_1 <= 5'h05;  // n (S 的近�?
                    digit_0 <= 5'h10;  // P
                end

                `GEN_RANDOM: begin
                    
                    digit_3 <= 5'h01;  // I
                    digit_2 <= 5'h05;  // n
                    digit_1 <= 5'h10;  // P
                    digit_0 <= 5'h11;  // t
                end

                `ERROR: begin
                    // ERROR״̬��ʾ�̶���"Err0"��������ά�ȳ�����Χʱ��ͬ��
                    // ������ʲô��������ά�ȴ������ݴ�������ά�Ȳ�ƥ�䣩������ʾ��ͬ����Ϣ
                    digit_3 <= 5'h0E;  // E
                    digit_2 <= 5'h13;  // r
                    digit_1 <= 5'h13;  // r
                    digit_0 <= 5'h00;  // 0����ʾ����
                end

                `BONUS: begin 
                    // ��BONUS״̬����ʾʱ����������cycles��
                    // ��ȡÿ��ʮ����λ��digit_3��ǧλ��digit_2�ǰ�λ��digit_1��ʮλ��digit_0�Ǹ�λ
                    // ������ʾ��ΧΪ0-9999��4λ���֣��������������ʾ9999
                    if (cycles > 32'd9999) begin
                        digit_3 <= 4'd9;
                        digit_2 <= 4'd9;
                        digit_1 <= 4'd9;
                        digit_0 <= 4'd9;
                    end else begin
                        digit_3 <= (cycles / 32'd1000) % 10;
                        digit_2 <= (cycles / 32'd100) % 10;
                        digit_1 <= (cycles / 32'd10) % 10;
                        digit_0 <= cycles % 10;
                    end
                end

                `OUTPUT_RES: begin
                    digit_3 <= 5'h00;  // o
                    digit_2 <= 5'h01;  // U
                    digit_1 <= 5'h11;  // t
                    digit_0 <= 5'h10;  // P
                end


                default: begin
                    digit_3 <= 5'h0F;
                    digit_2 <= 5'h0F;
                    digit_1 <= 5'h0F;
                    digit_0 <= 5'h0F;
                end
            endcase
        end
    end

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            led <= 8'b0;
        end
        else begin
            led <= 8'b0; 
            
            // ����LED���ȼ��������⵽����������ERROR״̬������led[7]
            if (error_led || (state == `ERROR)) begin
                if (state == `ERROR) 
                    led[7] <= refresh_cnt[19];  // ERROR״̬ʱ��˸
                else
                    led[7] <= 1'b1;  // �������ʱ������������
            end
            // ������ڴ���״̬�������״̬��ʾ��Ӧ��LED
            else begin
                case (state)
                    `IDLE:      led[0] <= 1'b1;
                    `INPUT_DIM: led[1] <= 1'b1;
                    `INPUT_DATA:led[2] <= 1'b1;
                    `FILL_ZEROS:led[2] <= 1'b1;
                    `COMPUTE:   led[3] <= 1'b1;
                    `BONUS:     led[4] <= 1'b1;
                    `OUTPUT_RES:led[5] <= 1'b1;
                    `DISPLAY_MODE: led[6] <= 1'b1;
                    `GEN_RANDOM: led[6] <= 1'b1;
                    default:    led <= 8'b0;
                endcase
            end
        end
    end

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            scan_cnt <= 2'd0;
            refresh_cnt <= 20'd0;
        end
        else begin
            refresh_cnt <= refresh_cnt + 1;
            if (refresh_cnt >= 20'd200_000) begin 
                refresh_cnt <= 0;
                scan_cnt <= scan_cnt + 1;
            end
        end
    end

    
    always @(*) begin
        an = 4'b0000;
        current_digit = 5'h00;

        case (scan_cnt)
            2'd0: begin
                an = 4'b0001;
                current_digit = digit_0;
            end
            2'd1: begin
                an = 4'b0010;
                current_digit = digit_1;
            end
            2'd2: begin
                an = 4'b0100;
                current_digit = digit_2;
            end
            2'd3: begin
                an = 4'b1000;
                current_digit = digit_3;
            end
            default: begin
                an = 4'b0000;
                current_digit = 5'h00;
            end
        endcase
    end

    
    always @(*) begin
        case (current_digit)
            5'h00: seg = 8'h3F; 
            5'h01: seg = 8'h06; 
            5'h02: seg = 8'h5B;
            5'h03: seg = 8'h4F;
            5'h04: seg = 8'h66;
            5'h05: seg = 8'h6D;
            5'h06: seg = 8'h7D;
            5'h07: seg = 8'h07;
            5'h08: seg = 8'h7F;
            5'h09: seg = 8'h6F;

            5'h0A: seg = 8'h77; //A
            5'h0B: seg = 8'h7C; //b
            5'h0C: seg = 8'h39; //C
            5'h0D: seg = 8'h5E; //d
            5'h0E: seg = 8'h79; //E
            5'h0F: seg = 8'h71; //F
            5'h10: seg = 8'h73; //P
            5'h11: seg = 8'h78; //t
            5'h12: seg = 8'h38; //L
            5'h13: seg = 8'h50; //r
            5'h14: seg = 8'h78; //T (same as t)
            5'h15: seg = 8'h1E; //J

            default: seg = 8'h00; //default默认全灭
        endcase
    end

endmodule
