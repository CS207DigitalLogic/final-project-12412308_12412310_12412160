`ifndef PARAMETERS_VH
`define PARAMETERS_VH


`define IDLE 0
`define INPUT_DIM 1
`define INPUT_DATA 2
`define FILL_ZEROS 7
`define COMPUTE 3
`define OUTPUT_RES 4
`define ERROR 5
`define BONUS 6
`define GEN_RANDOM 8
`define DISPLAY_MODE 9


// ASCII �?
`define ASCII_SPACE 8'h20
`define ASCII_NEWLINE 8'h0A
`define ASCII_CR 8'h0D
`define ASCII_MINUS 8'h2D
`define ASCII_0 8'h30
`define ASCII_9 8'h39
`define ASCII_E 8'h45  // 'E'
`define ASCII_R 8'h52  // 'R'
`define ASCII_O 8'h4F  // 'O'


`define MAX_ROWS 5
`define MAX_COLS 5
`define BIT_PERIOD 16'd867

`endif