`include "parameters.vh"

module input_image_rom(
    input clk,
    input [3:0] x,
    input [3:0] y,
    output reg [3:0] data_out
);

    reg [3:0] rom [0:119];

    initial begin 
        rom[0] = 4'd3;  rom[1] = 4'd7;  rom[2] = 4'd2;  rom[3] = 4'd9;  
        rom[4] = 4'd0;  rom[5] = 4'd5;  rom[6] = 4'd1;  rom[7] = 4'd8;  
        rom[8] = 4'd4;  rom[9] = 4'd6;  rom[10] = 4'd3; rom[11] = 4'd2;

        rom[12] = 4'd8; rom[13] = 4'd1; rom[14] = 4'd6; rom[15] = 4'd4; 
    rom[16] = 4'd7; rom[17] = 4'd3; rom[18] = 4'd9; rom[19] = 4'd0; 
    rom[20] = 4'd5; rom[21] = 4'd2; rom[22] = 4'd8; rom[23] = 4'd1; 

    
    rom[24] = 4'd4; rom[25] = 4'd9; rom[26] = 4'd0; rom[27] = 4'd2; 
    rom[28] = 4'd6; rom[29] = 4'd8; rom[30] = 4'd3; rom[31] = 4'd5; 
    rom[32] = 4'd7; rom[33] = 4'd1; rom[34] = 4'd4; rom[35] = 4'd9; 

    
    rom[36] = 4'd7; rom[37] = 4'd3; rom[38] = 4'd8; rom[39] = 4'd5; 
    rom[40] = 4'd1; rom[41] = 4'd4; rom[42] = 4'd9; rom[43] = 4'd2; 
    rom[44] = 4'd0; rom[45] = 4'd6; rom[46] = 4'd7; rom[47] = 4'd3; 

    
    rom[48] = 4'd2; rom[49] = 4'd6; rom[50] = 4'd4; rom[51] = 4'd0; 
    rom[52] = 4'd8; rom[53] = 4'd7; rom[54] = 4'd5; rom[55] = 4'd3; 
    rom[56] = 4'd1; rom[57] = 4'd9; rom[58] = 4'd2; rom[59] = 4'd4; 

    
    rom[60] = 4'd9; rom[61] = 4'd0; rom[62] = 4'd7; rom[63] = 4'd3; 
    rom[64] = 4'd5; rom[65] = 4'd2; rom[66] = 4'd8; rom[67] = 4'd6; 
    rom[68] = 4'd4; rom[69] = 4'd1; rom[70] = 4'd9; rom[71] = 4'd0; 

    
    rom[72] = 4'd5; rom[73] = 4'd8; rom[74] = 4'd1; rom[75] = 4'd6; 
    rom[76] = 4'd4; rom[77] = 4'd9; rom[78] = 4'd2; rom[79] = 4'd7; 
    rom[80] = 4'd3; rom[81] = 4'd0; rom[82] = 4'd5; rom[83] = 4'd8; 

    
    rom[84] = 4'd1; rom[85] = 4'd4; rom[86] = 4'd9; rom[87] = 4'd2; 
    rom[88] = 4'd7; rom[89] = 4'd0; rom[90] = 4'd6; rom[91] = 4'd8; 
    rom[92] = 4'd5; rom[93] = 4'd3; rom[94] = 4'd1; rom[95] = 4'd4; 

    
    rom[96] = 4'd6;  rom[97] = 4'd2;  rom[98] = 4'd5;  rom[99] = 4'd8;  
    rom[100]= 4'd3;  rom[101]= 4'd1;  rom[102]= 4'd7;  rom[103]= 4'd4; 
    rom[104]= 4'd9;  rom[105]= 4'd0;  rom[106]= 4'd6;  rom[107]= 4'd2; 

    
    rom[108]= 4'd0;  rom[109]= 4'd7;  rom[110]= 4'd3;  rom[111]= 4'd9; 
    rom[112]= 4'd5;  rom[113]= 4'd6;  rom[114]= 4'd4;  rom[115]= 4'd1; 
    rom[116]= 4'd8;  rom[117]= 4'd2;  rom[118]= 4'd0;  rom[119]= 4'd7; 
end


wire [6:0] addr; 

assign addr = x*12+y; 

always @(*) begin 
    data_out = rom[addr]; 
end 

endmodule
